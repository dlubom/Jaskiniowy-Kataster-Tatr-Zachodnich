++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
 A B I S S O  v5.0�
 Vypocet (a vyrovnanie) polyg�nov�ho merania jaskyne : OBC_VYV.SS
 
                                              DATE :  13- 8-2003/11:58:39
                                              SoftShip/Abisso PPP(C) 1996
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++

 N�zov syst�mu:  Jaskyna OBCASNA VYVIERACKA, Cervene vrchy

 Lokalita     :  Rozpadly grun, Cervene vrchy
 Zameral(i)   :  viacer�, skupina SSS Ruzomberok
 D�tum        :  13.8.1979

 TAH POLYGONU od bodu -1�>2 po bod 20 � 20 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   -1    72.00    53.00   118.00     0.00     0.00   1435.00    Pripojny bod
    2    72.23    53.18   116.00     2.02     0.30   1433.00  
    3    69.54    53.66   114.94     4.95     3.03   1431.94           
    4    56.94    54.09   114.88    17.56    15.64   1431.88  HLADINA I.SIFON
    5    49.20    56.10   112.81    25.82    23.63   1429.81  I.SIFON
    6    38.20    50.97   114.84    38.12    35.76   1431.84  SIEN I.-II.SIF.
    7    27.01    52.24   114.19    49.40    47.03   1431.19           
    8    15.41    52.24   113.99    61.01    58.63   1430.99           
    9     8.61    53.69   112.34    68.15    65.58   1429.34  II.SIFON
   10    -1.11    53.69   113.36    77.92    75.30   1430.36           
   11   -13.83    50.27   115.05    91.20    88.47   1432.05           
   12   -23.94    49.39   116.84   101.51    98.63   1433.84           
   13   -23.95    49.39   133.89   118.56    98.63   1450.89           
   14   -32.56    47.56   135.91   127.59   107.43   1452.91  SIEN OBJAVITEL.
   15   -32.50    45.85   132.62   131.30   109.14   1449.62  UZINA K JAZERU
   16   -38.91    45.73   130.16   138.17   115.55   1447.16           
   17   -42.84    51.15   128.17   145.15   122.25   1445.17  JAZERO 30cm POD
   18   -49.46    54.66   128.17   152.64   129.74   1445.17  KANAL
   19   -53.94    60.83   129.45   160.37   137.36   1446.45           
   20   -63.17    65.95   127.72   171.07   147.92   1444.72           

 Prevysenie  23.56  m b. imax=    14 a imin=     9, dlzka   171.07  m
________________________________________________________________________

 TAH POLYGONU od bodu 14�>21 po bod 22 � 22 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   14   -32.56    47.56   135.91     0.00     0.00   1452.91  SIEN OBJAVITEL.
   21   -27.69    42.86   133.71     7.11     6.76   1450.71  SIEN OBJAVITEL.
   22   -25.83    41.30   133.52     9.55     9.19   1450.52  PIESOCNA CHODB.

 Prevysenie   2.39  m b. imax=    14 a imin=    22, dlzka     9.55  m
________________________________________________________________________

 TAH POLYGONU od bodu 14�>23 po bod 23 � 23 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   14   -32.56    47.56   135.91     0.00     0.00   1452.91  SIEN OBJAVITEL.
   23   -27.33    46.06   135.19     5.48     5.43   1452.19  S.O.

 Prevysenie   0.72  m b. imax=    14 a imin=    23, dlzka     5.48  m
________________________________________________________________________

 TAH POLYGONU od bodu 14�>24 po bod 24 � 24 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   14   -32.56    47.56   135.91     0.00     0.00   1452.91  SIEN OBJAVITEL.
   24   -29.37    51.64   134.62     5.34     5.18   1451.62  S.O.

 Prevysenie   1.29  m b. imax=    14 a imin=    24, dlzka     5.34  m
________________________________________________________________________

 TAH POLYGONU od bodu 14�>25 po bod 25 � 25 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   14   -32.56    47.56   135.91     0.00     0.00   1452.91  SIEN OBJAVITEL.
   25   -33.60    50.29   134.79     3.13     2.92   1451.79  S.O.

 Prevysenie   1.12  m b. imax=    14 a imin=    25, dlzka     3.13  m
________________________________________________________________________

 TAH POLYGONU od bodu 14�>26 po bod 27 � 27 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   14   -32.56    47.56   135.91     0.00     0.00   1452.91  SIEN OBJAVITEL.
   26   -26.60    50.72   144.69    11.07     6.74   1461.69  Horne vetvy
   27   -20.75    49.04   145.93    17.29    12.83   1462.93           

 Prevysenie  10.02  m b. imax=    27 a imin=    14, dlzka    17.29  m
________________________________________________________________________

 TAH POLYGONU od bodu 26�>28 po bod 28 � 28 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   26   -26.60    50.72   144.69     0.00     0.00   1461.69  Horne vetvy
   28   -23.06    54.40   147.46     5.81     5.11   1464.46  VODOPAD

 Prevysenie   2.77  m b. imax=    28 a imin=    26, dlzka     5.81  m
________________________________________________________________________

 TAH POLYGONU od bodu 26�>29 po bod 31 � 31 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   26   -26.60    50.72   144.69     0.00     0.00   1461.69  Horne vetvy
   29   -29.76    55.23   144.59     5.50     5.50   1461.59           
   30   -26.65    59.07   148.70    11.92    10.44   1465.70           
   31   -22.59    59.49   151.15    16.68    14.52   1468.15  SPOJENIE K B_27

 Prevysenie   6.55  m b. imax=    31 a imin=    29, dlzka    16.68  m
________________________________________________________________________

 TAH POLYGONU od bodu 30�>32 po bod 34 � 34 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   30   -26.65    59.07   148.70     0.00     0.00   1465.70           
   32   -25.69    61.85   149.92     3.19     2.95   1466.92           
   33   -30.41    66.91   152.12    10.45     9.87   1469.12           
   34   -27.45    66.28   156.37    15.67    12.90   1473.37  PRITOKOVY KOMIN

 Prevysenie   7.67  m b. imax=    34 a imin=    30, dlzka    15.67  m
________________________________________________________________________

 TAH POLYGONU od bodu 20�>35 po bod 40 � 40 (OTVORENY)

    #      x        y        z       dl        r     n.m.v.
    -      m        m        m        m        m         m
   20   -63.17    65.95   127.72     0.00     0.00   1444.72           
   35   -72.03    69.17   124.57     9.94     9.43   1441.57  III.SIFON
   36   -73.94    66.12   124.98    13.56    13.02   1441.98           
   37   -78.83    63.30   130.06    21.16    18.67   1447.06  REBRIK
   38   -81.06    61.42   130.01    24.08    21.59   1447.01  
   39   -86.15    68.97   122.64    35.79    30.69   1439.64  IV.SIFON-PLAZ
   40   -84.80    74.41   119.89    42.04    36.30   1436.89  24cm nad hladin.

 Prevysenie  10.17  m b. imax=    37 a imin=    40, dlzka    42.04  m
________________________________________________________________________


 DENIVELACIA SYSTEMU      44.02  m,  b.iMAX=    34, n.m.v.:  1473.37  m
                                     b.iMIN=     9, n.m.v.:  1429.34  m

 V KVADRI S ROZMERMI X:   158.39 m x Y:    33.11 m x Z:    44.02 m
 POCET VETIEV MERANIA :    10, v tom      0 vyrovnanych

 CELKOVA DLZKA SYSTEMU    292.06  m NA     40 BODOCH
 & 
